package Testing;

endpackage
