package Endian;

import Vector::*;
import StmtFSM::*;

typedef union tagged {
    void Unused00;
    Bit#(64) Bit64_01;
    void Unused02;
    void Unused03;
    void Unused04;
    void Unused05;
    void Unused06;
    void Unused07;
    void Unused08;
    void Unused09;
    void Unused0A;
    void Unused0B;
    void Unused0C;
    void Unused0D;
    void Unused0E;
    void Unused0F;
    void Unused10;
    void Unused11;
    void Unused12;
    void Unused13;
    void Unused14;
    void Unused15;
    void Unused16;
    void Unused17;
    void Unused18;
    void Unused19;
    void Unused1A;
    void Unused1B;
    void Unused1C;
    void Unused1D;
    void Unused1E;
    void Unused1F;
    void Unused20;
    void Unused21;
    void Unused22;
    void Unused23;
    void Unused24;
    void Unused25;
    void Unused26;
    void Unused27;
    void Unused28;
    void Unused29;
    void Unused2A;
    void Unused2B;
    void Unused2C;
    void Unused2D;
    void Unused2E;
    void Unused2F;
    void Unused30;
    void Unused31;
    void Unused32;
    void Unused33;
    void Unused34;
    void Unused35;
    void Unused36;
    void Unused37;
    void Unused38;
    void Unused39;
    void Unused3A;
    void Unused3B;
    void Unused3C;
    void Unused3D;
    void Unused3E;
    void Unused3F;
    void Unused40;
    void Unused41;
    void Unused42;
    void Unused43;
    void Unused44;
    void Unused45;
    void Unused46;
    void Unused47;
    void Unused48;
    void Unused49;
    void Unused4A;
    void Unused4B;
    void Unused4C;
    void Unused4D;
    void Unused4E;
    void Unused4F;
    void Unused50;
    void Unused51;
    void Unused52;
    void Unused53;
    void Unused54;
    void Unused55;
    void Unused56;
    void Unused57;
    void Unused58;
    void Unused59;
    void Unused5A;
    void Unused5B;
    void Unused5C;
    void Unused5D;
    void Unused5E;
    void Unused5F;
    void Unused60;
    void Unused61;
    void Unused62;
    void Unused63;
    void Unused64;
    void Unused65;
    void Unused66;
    void Unused67;
    void Unused68;
    void Unused69;
    void Unused6A;
    void Unused6B;
    void Unused6C;
    void Unused6D;
    void Unused6E;
    void Unused6F;
    void Unused70;
    void Unused71;
    void Unused72;
    void Unused73;
    void Unused74;
    void Unused75;
    void Unused76;
    void Unused77;
    void Unused78;
    void Unused79;
    void Unused7A;
    void Unused7B;
    void Unused7C;
    void Unused7D;
    void Unused7E;
    void Unused7F;
    void Unused80;
    void Unused81;
    void Unused82;
    void Unused83;
    void Unused84;
    void Unused85;
    void Unused86;
    void Unused87;
    void Unused88;
    void Unused89;
    void Unused8A;
    void Unused8B;
    void Unused8C;
    void Unused8D;
    void Unused8E;
    void Unused8F;
    void Unused90;
    void Unused91;
    void Unused92;
    void Unused93;
    void Unused94;
    void Unused95;
    void Unused96;
    void Unused97;
    void Unused98;
    void Unused99;
    void Unused9A;
    void Unused9B;
    void Unused9C;
    void Unused9D;
    void Unused9E;
    void Unused9F;
    void UnusedA0;
    void UnusedA1;
    void UnusedA2;
    void UnusedA3;
    void UnusedA4;
    void UnusedA5;
    void UnusedA6;
    void UnusedA7;
    void UnusedA8;
    void UnusedA9;
    void UnusedAA;
    void UnusedAB;
    void UnusedAC;
    void UnusedAD;
    void UnusedAE;
    void UnusedAF;
    void UnusedB0;
    void UnusedB1;
    void UnusedB2;
    void UnusedB3;
    void UnusedB4;
    void UnusedB5;
    void UnusedB6;
    void UnusedB7;
    void UnusedB8;
    void UnusedB9;
    void UnusedBA;
    void UnusedBB;
    void UnusedBC;
    void UnusedBD;
    void UnusedBE;
    void UnusedBF;
    void UnusedC0;
    void UnusedC1;
    void UnusedC2;
    void UnusedC3;
    void UnusedC4;
    void UnusedC5;
    void UnusedC6;
    void UnusedC7;
    void UnusedC8;
    void UnusedC9;
    void UnusedCA;
    void UnusedCB;
    void UnusedCC;
    void UnusedCD;
    void UnusedCE;
    void UnusedCF;
    void UnusedD0;
    void UnusedD1;
    void UnusedD2;
    void UnusedD3;
    void UnusedD4;
    void UnusedD5;
    void UnusedD6;
    void UnusedD7;
    void UnusedD8;
    void UnusedD9;
    void UnusedDA;
    void UnusedDB;
    void UnusedDC;
    void UnusedDD;
    void UnusedDE;
    void UnusedDF;
    void UnusedE0;
    void UnusedE1;
    void UnusedE2;
    void UnusedE3;
    void UnusedE4;
    void UnusedE5;
    void UnusedE6;
    void UnusedE7;
    void UnusedE8;
    void UnusedE9;
    void UnusedEA;
    void UnusedEB;
    void UnusedEC;
    void UnusedED;
    void UnusedEE;
    void UnusedEF;
    void UnusedF0;
    void UnusedF1;
    void UnusedF2;
    void UnusedF3;
    void UnusedF4;
    void UnusedF5;
    void UnusedF6;
    void UnusedF7;
    void UnusedF8;
    void UnusedF9;
    Bit#(32) Bit32_FA;
    void UnusedFB;
    void UnusedFC;
    void UnusedFD;
    void UnusedFE;
    void UnusedFF;
} Union8b deriving(Eq,FShow,Bits);

typedef struct {
    Bit#(64) a64;
    Bit#(32) b32;
    Bit#(32) c32;
} Foo deriving (Bits);


module mkTB_PrintEndian();

    Bit#(128) b = 128'h000102030405060708090a0b0c0d0e0f;

    Stmt masterstmt = seq
        $display("Bluespec packing conventions");
        $display("============================");
        $display;

        $display("  UnusedFC packs to: %018X",pack(tagged UnusedFC));
        $display("  Unused00 packs to: %018X",pack(tagged UnusedFC));
        $display("  Bit64_01 packs to: %018X",pack(tagged Bit64_01 64'hdeadbeef01234567));
        $display("  Bit32_FA packs to: %018X",pack(tagged Bit32_FA 32'h01234567));
        $display("  Unions pack with the tag at the MSB, [Pmax:P] padding and the payload at [P-1:0]");
        $display;
        action
            Union8b u = tagged Bit32_FA 32'h11111111;
            $display("  Bit32_FA with all 1's: fshow='",fshow(u),"'");
            $display("  Bit32_FA accessed by .Bit64_01: ",fshow(u.Bit64_01));
            $display("  Bit32_FA accessed by .Bit32_FA: ",fshow(u.Bit32_FA));
            $display("  Accessing by the wrong tag returns X");
        endaction
        $display;

        $display("Maybe#(Bit#(32))");
        $display("  32b tagged invalid packs to: %09X",pack(Maybe#(Bit#(32))'(tagged Invalid)));
        $display("  32b tagged valid   packs to: %09X",pack(Maybe#(Bit#(32))'(tagged Valid 32'h01234567)));
        $display("  Maybe#(t) is stored with a valid bit, followed by the data");
        $display;

        $display("b = %032X",b);
        action
            Vector#(2,Bit#(64)) p = unpack(b);
            $display("  As two 64b vectors: p[1]=%016X",p[1]);
            $display("                      p[0]=%016X",p[0]);
            $display("  Vectors are stored with highest index at MSB");
            $display;
        endaction

        action
            Foo t = unpack(b);
            $display("  As struct: a64=%16X b32=%8X c32=%8X",t.a64,t.b32,t.c32);
            $display("  Structs are stored with first element at MSB");
            $display;
        endaction

        action
            Tuple2#(Bit#(64),Bit#(64)) t = unpack(b);
            $display("  As Tuple2#(Bit#(64),Bit#(64)): first=%016X, second=%016X",tpl_1(t),tpl_2(t));
            $display("  Tuples are stored with the first element at MSB");
            $display;
        endaction

    endseq;

    mkAutoFSM(masterstmt);

endmodule

endpackage
